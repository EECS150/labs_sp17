module structural_adder (
    input [7:0] a,
    input [7:0] b,
    output [8:0] sum
);
    // Remove this line once you have implemented the structural adder
    assign sum = 9'd0;

endmodule
