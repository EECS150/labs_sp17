module rotary_decoder (
    input clk,
    input rst,
    input rotary_A,
    input rotary_B,
    output rotary_event,
    output rotary_left
);

    // Create your rotary decoder circuit here
    // This module takes in rotary_A and rotary_B which are the A and B signals synchronized to clk

    // Remove these lines after implementing your rotary decoder
    assign rotary_event = 0;
    assign rotary_left = 0;
endmodule
